-------------------------------------------------------------------------------
--
-- Title       : rs_in
-- Design      : rs_in
-- Author      : 
-- Company     : 
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_unsigned.all;--!!!!!!!!!!!!!!!!!! ������ �������� �� ��� �������! ��� ����� ��� �������� ����   cnt<= cnt+ '1';

entity rs_in is	  
	port(
	clk			: in std_logic;  --100Mhz
	reset		: in std_logic;  -- 1 - reset
	uart_in		: in std_logic;
	data_out	: out std_logic_vector(7 downto 0);
	data_rdy	: out std_logic
	);
end rs_in;			



architecture rs_in of rs_in is 
constant half_start_bit	: std_logic_vector(15 downto 0):=x"01B2"; -- ��� ��� ������. ������ �������� ����� ��������� � ����������� �� ����������� ������ UART � clk.
constant length_bit	: std_logic_vector(15 downto 0):=x"0361"; -- ��� ��� ������. ������ �������� ����� ��������� � ����������� �� ����������� ������ UART � clk.
constant uart_length	: std_logic_vector(3 downto 0):=x"7"; -- ����� ������� UART � �����
-- ���� �������� ��� ������� ��������, ������ x"2F6", �� ����� 16 �������� ��� ������� �������� �������� ������. 
-- ���������� ����� ������ 10 ��� 
signal cnt0			: std_logic_vector(15 downto 0); -- ������� ������� ���������� ����  
signal cnt1			: std_logic_vector(15 downto 0); --������� �������� ��������� ����� ������ 
signal cnt_bits		: std_logic_vector(7 downto 0);  --������� ����������� ���

signal st_main		: std_logic_vector(1 downto 0):="00";		--������, ������������ ������ ��������� ��������. ����� �� ����� 4 ���������
signal shift_reg	: std_logic_vector(7 downto 0);

-- ������� ������� ��������
function reverse(X : in std_logic_vector) return std_logic_vector is
variable ret : std_logic_vector(X'range);
begin
    for i in X'range loop
        ret(i) := X(X'left - i);
    end loop;
   return ret;
end function;

begin
	
pr_main: process(clk)
	
begin  
	if(rising_edge(clk))then --��� ��������� ������ ������� if, ���� ���� ����������
		if(reset = '1')then  -- ���������� ��������� ������� � ���������� �������� �� ������
			st_main	<= "00";  --������, ������������ ������ ��������� ��������. ����� �� ����� 4 ���������
			data_rdy	<= '0';	-- ������ ��������� ������ ���������� �������� ������ �� ������ ��������. ����� ����� �������� ����������� ����������� �����. ������� ���������� ���� ������  
			cnt0	<= (others=>'0');	 
			data_out	<= (others=>'0');
		else   
			case st_main is 
			when "00"=>	  --��������� ���������. ���� ��������� ���
				if(	uart_in = '0')then --���� ������ ��������� ���, �������� ������� �������� ����� ����� ���������� ����, ���� ��������� ����������� ������ � ��������
					-- ���� ����� �� �������, �� � ���� ������������� ���������� ����� � ����� ������� ���������� �� ������ ���� � ������ � 
					-- ������� ������������ ��������� ����. �������� ��� ��������� �� ������� ��������� UART
					cnt0<= cnt0+ '1';  
				else
					cnt0	<= (others=>'0'); --���� ��� ������ uart_in = 0, �� �� ��� �������� uart_in � 1 ������� �������. ������ ������������ ����� ���������� ��-�� �������������  ����������� ����������
					--� ���. ��������, ���������� ����� ����������, � �� ������ ����� �����. ������ ������ ������������ �� ��������.																		 		
				end if;
				if( cnt0 = half_start_bit)then --���� �� ��������� �� ������� ��������, �� ��������� ���������� ���������� ���� 
					st_main	<= "01";	 --��������� � ��������� ����������� �������� ������� ������������ ����
					--cnt0 <=(others=>'0'); -- ����� �������� ������� ���������� ����
				end if;	 
				cnt1		<= (others=> '0'); --����� �������� ��� �������� ��������� ����� ������
				cnt_bits	<= (others=> '0'); --����� �������� �������
				--shift_reg  	<= (others=> '0'); --����� ���������� ��������
				data_rdy	<= '0';					
			when "01"=>	--����������� �������� ������� ������������ ����
				if( cnt1 = length_bit)then --���� �� ��������� �� ������� ��������, �� ������������� �� ������ ���� � ������ 
					st_main	<= "10";	 --��������� � ��������� ������������� ������� uart
				end if;	
				cnt1<= cnt1+ '1';  
				cnt0 <=(others=>'0'); -- ����� �������� ������� ���������� ����
			when "10"=>	--������������� ������� uart
				if(cnt_bits = uart_length)then 	  
					st_main	<= "11";-- ���� ������� ��� 8 ���, �� ��������� � ��������� ���������, � ������� ������� ������ ����������		
				else   
					st_main	<= "01";-- ��� 8 ��� ��� �� �������, ���� ��������� ��������� ���
				end if;
				cnt1		<= (others=> '0'); --����� �������� ��� �������� ��������� ����� ������
				shift_reg	<= shift_reg(6 downto 0) & uart_in; -- �������� ������ �����. ���������� ��������� ������� ��������� ������	 
				cnt_bits <= cnt_bits + '1'; -- ��������� ��� ������, ������ ����������� ������� �������� ���
			when "11"=>	  -- ������� ������� ���, ��������� ��������� ������� ������
				if(uart_in = '1')then  -- ���� �� ���� ������ �������� ���, �� ��������� � ��������� ��������� ��� ������ ���������� ���������� ����	
					st_main		<= "00"; -- 	
					data_rdy	<= '1';	
				else
					--����� �� ��������, ���� ���� ���� �� ����� ���.
				end if;
				data_out	<= reverse(shift_reg);--������ ������������������ ��� ��� �������� MSB  � LSB
				--data_out	<= shift_reg;
				--data_rdy	<= '1';			
			
			when others=> null;
			end case;
		end if;
		
				  
		
	end if;
	
end process;



end rs_in;
